library IEEE;
use IEEE.std_logic_1164.ALL;

entity total_tb is
end total_tb;

