library IEEE;
use IEEE.std_logic_1164.ALL;

entity chip_tb is
end chip_tb;

