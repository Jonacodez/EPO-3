library IEEE;
use IEEE.std_logic_1164.ALL;

entity detect_input is
port(   
	KEY0 : in std_logic;
	KEY1 : in std_logic;
	KEY2 : in std_logic;
	KEY3 : in std_logic;
	input_s : out std_logic
     );
end entity;


